module scoreboard_4_bit #(parameter DATA_WIDTH = 4, GOLDEN_WIDTH = 8, INPUT_WIDTH = 11);

    reg [INPUT_WIDTH-1:0] input_data [0:2047]; 
    reg [GOLDEN_WIDTH-1:0] golden [0:2047];  
    reg signed [DATA_WIDTH-1:0] a, b; 
    reg clk, reset;  
    reg [2:0] op;                        
    wire signed [GOLDEN_WIDTH-1:0] result;  
    reg signed [GOLDEN_WIDTH-1:0] expected;  
    integer i, mismatch_count, right_add, right_sub, right_mul, right_div;   
               

    ALU_standard_caculator_n_bit #(DATA_WIDTH) alu (
        .a(a),
        .b(b),
        .clk(clk),
        .rst(reset),
        .op(op),
        .result(result)
    );

    // initial clk = 1;
    always #5 clk = ~clk; 

    initial begin
        mismatch_count = 0;
        right_add = 0; right_sub = 0; right_mul = 0; right_div = 0;
        clk = 0;
        reset = 1; 

        $readmemb("E:/Code/Learn/Verilog/Homework/ALU n bit/ALU standard/input_signed.txt", input_data);
        $display("%b", input_data[0][INPUT_WIDTH-1:INPUT_WIDTH-DATA_WIDTH]);
        $readmemb("E:/Code/Learn/Verilog/Homework/ALU n bit/ALU standard/golden.txt", golden);

        #10 reset = 0;
        // #10;
        for (i = 0; i < 2048; i = i + 1) begin
            // reset = 1;
            a = input_data[i][INPUT_WIDTH-1:INPUT_WIDTH-DATA_WIDTH];
            b = input_data[i][INPUT_WIDTH-1-DATA_WIDTH:DATA_WIDTH-1];
            op = input_data[i][DATA_WIDTH-2:0];
            expected = golden[i];
            reset = 1;
            #5; reset = 0; 
            #(DATA_WIDTH*10+20-5);
            
            if (result !== expected) begin
                $display("Mismatch at index %0d: a = %d, b = %d, op = %d, Output = %d, Expected = %d",
                         i, a, b, op, result, expected);
                mismatch_count = mismatch_count + 1;
            end else begin
                $display("Match at index %0d: a = %d, b = %d, op = %d, Output = %d, Expected = %d",
                         i, a, b, op, result, expected);
                case (op)
                    3'b000: right_add = right_add + 1;
                    3'b001: right_sub = right_sub + 1;
                    3'b010: right_mul = right_mul + 1;
                    3'b011: right_div = right_div + 1; 
                    default: right_add = right_add;
                endcase
            end
        end

        if (mismatch_count == 0) begin
            $display("All outputs match the golden file. Multiplier is correct.");
            $display("

@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@..@@@@@@@@@@@@@@@@@ :@@@@@@@@@@@@@@@@@@:.@@@@@@@@@@@@@@@@@@..@@@@@@@@@@@@@@@@@ .@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@::@@@@@@@@@@@@@@@@@.: @@@@@@@@@@@@@@@@@..@@@@@@@@@@@@@@@@@ ::@@@@@@@@@@@@@@@@@:: @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.::.@@@@@@@@@@@@@@@@::.@@@@@@@@@@@@@@@@ :: @@@@@@@@@@@@@@@@.::@@@@@@@@@@@@@@@@ ::.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@::::@@@@@@@@@@@@@@@@::: @@@@@@@@@@@@@@@ :: @@@@@@@@@@@@@@@ :::@@@@@@@@@@@@@@@@::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.:::::::::::::@@@@@ :::::::::::::@@@@@@::::::::::::::@@@@@@::::::::::::: @@@@@.:::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.::::::::::::.@@@@@ .::::::::::::@@@@@@::::::::::::::@@@@@@::::::::::::. @@@@@.:::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ :::::::::: @@@@@@@@::::::::::.@@@@@@@@ .::::::::: @@@@@@@@ ::::::::::@@@@@@@@ ::::::::::.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ .::::::: @@@@@@@@@@ ::::::::@@@@@@@@@@ ::::::::=@@@@@@@@@@:::::::::@@@@@@@@@@@.::::::: @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.::::::.@@@@@@@@@@@@::::::.@@@@@@@@@@@@@:::::: @@@@@@@@@@@@.::::::@@@@@@@@@@@@ ::::::.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@::::::::@@@@@@@@@@@@::::::: @@@@@@@@@@@ :::::: @@@@@@@@@@@@:::::::@@@@@@@@@@@@.:::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@::::::::@@@@@@@@@@@ ::: :::.@@@@@@@@@@@:::. :::@@@@@@@@@@@ ::: ::: @@@@@@@@@@@::::.:::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ::.@@.::@@@@@@@@@@@.::@@ :::@@@@@@@@@@ :::@@::: @@@@@@@@@@:::-@@.:.@@@@@@@@@@@::.@@ :: @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ .@@@@@ : @@@@@@@@@@: @@@@@. @@@@@@@@@@..@@@@@@..@@@@@@@@@@..@@@@@ :@@@@@@@@@@@: @@@@ . @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@.::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::@@@@@:::::::::::.@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@:::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::.@@@@.::::::::::: @@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@:::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::@@@@ :::::::::::.@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@ ::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::@@@@.::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@:::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::@@@@ :::::::::::: @@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@ :::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::.@@@ ::::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::: @@@.::::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::: @@ .:::::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.:::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::::: @ .:::::::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  ................................................:::::::::::. @@@@@......:::::::::::.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ :::::::::::.@@@@@@@@@@@@::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@...:.....:::::::::::::::::::::::::::::::::.  .:::::::::::@@@@@@@@@@@@.:::::::::::.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ .::::::::::::::::::::::::::::::::::::::::: :::::::::::: @@@@@@@@@@@ ::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@::::::::::::::::::::::::::::::::::::::::  ::::::::::::@@@@@@@@@@@@::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ::::::::::::::::::::::::::::::::::::::.@:::::::::::.@@@@@@@@@@@@ ::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ .:::::::::::::::::::::::::::::::::::@.:::::::::::@@@@@@@@@@@@ :::::::::::.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ..  .    ...      ....    . .. :@ :::::::::::.@@@@@@@@@@@@::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.............................:@ :::::::::::.@@@@@@@@@@@@.:::::::::::.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.:::::::::::::::::::::::::::: @::::::::::::@@@@@@@@@@@@.:::::::::::.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ::::::::::::::::::::::::::::@.:::::::::::.@@@@@@@@@@@@::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.::::::::::::::::::::::::::. ::::::::::::@@@@@@@@@@@@ :::::::::::.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.:::::::::::::::::::::::.@:::::::::::.@@@@@@@@@@@@:::::::::::: @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ::::::::::::::::::::::@ ::::::::::::@@@@@@@@@@@@.:::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.::::::::::: @@@@@@@@@@@@.::::::::::: @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.::::::::::::::::@@::::::::::::@@@@@@@@@@@@.:::::::::::.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ::::::::::::::::@.::::::::::: @@@@@@@@@@@@::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@:::::::::::::::: ::::::::::::@@@@@@@@@@@@.:::::::::::-@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ::::::::::::.@::::::::::::@@@@@@@@@@@@:::::::::::: @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ :::::::::::@ :::::::::::.@@@@@@@@@@@@::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@       @:::::::::::: @@@@@@@@@@@@:::::::::::: @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.:::::::::::@@@@@@@@@@@@.::::::::::: @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.::::::::::: @@@@@@@@@@@ ::::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.:::::::::::.@@@@@@@@@@@@.::::::::::: @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@::::::::::::@@@@@@@@@@@@ ::::::::::: @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@::::::::::: @@@@@@@@@@@@.::::::::::.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@:::::::::: @@@@@@@@@@@@@ ::::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@.:::::::::@@@@@@@@@@@@@@@::::::::: @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@:::::::: @@@@@@@@@@@@@@@ ::::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ ::::::.@@@@@@@@@@@@@@@@@.::::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@ :::::@@@@@@@@@@@@@@@@@@@ ::::@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@::: @@@@@@@@@@@@@@@@@@@@:::.@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@
            
            ");
            $display("ADD right is : %d / 256", right_add);
            $display("SUB right is : %d / 256", right_sub);
            $display("MUL right is : %d / 256", right_mul);
            $display("DIV right is : %d / 256", right_div);
        end else begin
            $display("Multiplier is incorrect. Total mismatches: %0d", mismatch_count);
            $display("ADD right is : %d / 256", right_add);
            $display("SUB right is : %d / 256", right_sub);
            $display("MUL right is : %d / 256", right_mul);
            $display("DIV right is : %d / 256", right_div);
            
        end

        $stop;
    end
endmodule
